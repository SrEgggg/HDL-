module XOR_gate_level(output Y, input A, B);
  xor(Y, A, B);  // Built-in XOR primitive
endmodule
