module OR_data_flow (output Y, input A, B, C);
	assign Y = A || B || C;
endmodule