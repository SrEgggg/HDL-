module XOR_data_flow(output Y, input A, B);
  // Dataflow modeling of XOR
  assign Y = A ^ B;
endmodule
