module XNOR_gate_level(output Y, input A, B);
  xnor(Y, A, B);  // Built-in XNOR primitive
endmodule
