module OR_gate_level (output Y, input A, B, C);
	or(Y, A, B, C);
endmodule