module NOR_2_data_flow(output Y,input A,B);
	assign Y = ~ (A | B);
endmodule;