module NAND_gate_level(output Y, input A, B);
  nand(Y, A, B); 
endmodule
